library verilog;
use verilog.vl_types.all;
entity lab1_5_vlg_vec_tst is
end lab1_5_vlg_vec_tst;
