library verilog;
use verilog.vl_types.all;
entity lab4_1_vlg_vec_tst is
end lab4_1_vlg_vec_tst;
