library verilog;
use verilog.vl_types.all;
entity lab1_1 is
    port(
        sw0             : in     vl_logic;
        sw1             : in     vl_logic;
        sw2             : in     vl_logic;
        led0            : out    vl_logic;
        led1            : out    vl_logic;
        led2            : out    vl_logic;
        led3            : out    vl_logic;
        led4            : out    vl_logic;
        led5            : out    vl_logic;
        led6            : out    vl_logic;
        led7            : out    vl_logic;
        led8            : out    vl_logic;
        led9            : out    vl_logic
    );
end lab1_1;
