library verilog;
use verilog.vl_types.all;
entity lab1_1_vlg_check_tst is
    port(
        led0            : in     vl_logic;
        led1            : in     vl_logic;
        led2            : in     vl_logic;
        led3            : in     vl_logic;
        led4            : in     vl_logic;
        led5            : in     vl_logic;
        led6            : in     vl_logic;
        led7            : in     vl_logic;
        led8            : in     vl_logic;
        led9            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab1_1_vlg_check_tst;
