module test

(input signed [7:0] a,
input real [7:0] b,
output [15:0] res);

assign res =  a*b;


endmodule 